library verilog;
use verilog.vl_types.all;
entity project5_vlg_vec_tst is
end project5_vlg_vec_tst;
