library verilog;
use verilog.vl_types.all;
entity project8_vlg_vec_tst is
end project8_vlg_vec_tst;
