library verilog;
use verilog.vl_types.all;
entity KS8_vlg_vec_tst is
end KS8_vlg_vec_tst;
