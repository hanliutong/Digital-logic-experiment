library verilog;
use verilog.vl_types.all;
entity project6 is
    port(
        a               : out    vl_logic;
        CLK             : in     vl_logic;
        reset           : in     vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic;
        ds1             : out    vl_logic;
        ds2             : out    vl_logic;
        RCO             : out    vl_logic
    );
end project6;
