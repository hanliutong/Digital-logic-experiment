library verilog;
use verilog.vl_types.all;
entity BCDplus_vlg_vec_tst is
end BCDplus_vlg_vec_tst;
