library verilog;
use verilog.vl_types.all;
entity test_vlg_check_tst is
    port(
        out_test        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end test_vlg_check_tst;
