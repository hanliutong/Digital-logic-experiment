library verilog;
use verilog.vl_types.all;
entity decoder2_3_vlg_vec_tst is
end decoder2_3_vlg_vec_tst;
