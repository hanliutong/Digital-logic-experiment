library verilog;
use verilog.vl_types.all;
entity project3_vlg_vec_tst is
end project3_vlg_vec_tst;
