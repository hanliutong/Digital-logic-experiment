library verilog;
use verilog.vl_types.all;
entity count_B32_vlg_vec_tst is
end count_B32_vlg_vec_tst;
