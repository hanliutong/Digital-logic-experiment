library verilog;
use verilog.vl_types.all;
entity Verilog1_vlg_check_tst is
    port(
        F_C             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Verilog1_vlg_check_tst;
