library verilog;
use verilog.vl_types.all;
entity project9_vlg_vec_tst is
end project9_vlg_vec_tst;
