library verilog;
use verilog.vl_types.all;
entity project9_vlg_check_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        DS1             : in     vl_logic;
        DS2             : in     vl_logic;
        DS3             : in     vl_logic;
        DS4             : in     vl_logic;
        DS5             : in     vl_logic;
        DS6             : in     vl_logic;
        DS7             : in     vl_logic;
        DS8             : in     vl_logic;
        E               : in     vl_logic;
        F               : in     vl_logic;
        G               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end project9_vlg_check_tst;
