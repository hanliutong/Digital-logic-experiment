library verilog;
use verilog.vl_types.all;
entity decoder2_4_vlg_vec_tst is
end decoder2_4_vlg_vec_tst;
