library verilog;
use verilog.vl_types.all;
entity motor_12_vlg_vec_tst is
end motor_12_vlg_vec_tst;
