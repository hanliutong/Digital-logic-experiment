library verilog;
use verilog.vl_types.all;
entity kbd_vlg_vec_tst is
end kbd_vlg_vec_tst;
