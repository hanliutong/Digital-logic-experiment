library verilog;
use verilog.vl_types.all;
entity Verilog1_vlg_vec_tst is
end Verilog1_vlg_vec_tst;
