library verilog;
use verilog.vl_types.all;
entity project4_vlg_vec_tst is
end project4_vlg_vec_tst;
