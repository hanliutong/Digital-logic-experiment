library verilog;
use verilog.vl_types.all;
entity floor_vlg_vec_tst is
end floor_vlg_vec_tst;
