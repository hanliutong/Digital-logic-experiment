library verilog;
use verilog.vl_types.all;
entity adder8_vlg_vec_tst is
end adder8_vlg_vec_tst;
