library verilog;
use verilog.vl_types.all;
entity register8_vlg_vec_tst is
end register8_vlg_vec_tst;
