module dot_matrix_ev(Fin_1up,Fin_2up,Fin_3up,Fin_2dn,Fin_3dn,Fin_4dn,Fin_1,Fin_2,Fin_3,Fin_4,drc,clk,row,col,door,c_floor,err);
input door,err;
input Fin_1up,Fin_2up,Fin_3up;
input Fin_2dn,Fin_3dn,Fin_4dn;
input Fin_1,Fin_2,Fin_3,Fin_4;
input [1:0]drc,c_floor;
input clk;
output reg [15:0] row;//行数据信号
output reg [3:0] col;//列扫描信号
reg clk1,clk2;
reg [1:0]cnt_d;
integer i,j;
reg [15:0]    r[0:99];
reg [7:0]    R[0:99];
initial 
   begin
     col=4'b1111; row=16'b0; 
	end
	
always @(posedge clk1)//字库
   begin
      R[0]=8'b0001_0000;R[1]=8'b0010_0000;R[2]=8'b0100_0000;
		R[3]=8'b1111_1111;R[4]=8'b0100_0000;R[5]=8'b0010_0000;
		R[6]=8'b0001_0000;R[7]=8'b0000_0000;//上箭头
		
		R[8]=8'b0000_1000;R[9]=8'b0000_0100;R[10]=8'b0000_0010;
		R[11]=8'b1111_1111;R[12]=8'b0000_0010;R[13]=8'b0000_0100;
		R[14]=8'b0000_1000;R[15]=8'b0000_0000;//下箭头

		R[16]=8'b0001_1000;//横杠
		
		R[17]=8'b0000_0000;R[18]=8'b0010_0010;R[19]=8'b0111_1110;
		R[20]=8'b0000_0010;R[21]=8'b0000_0000;R[22]=8'b0000_0000;
		R[23]=8'b0000_0000;R[24]=8'b0000_0000;//数字1
	
		R[25]=8'b0000_0000;R[26]=8'b0010_0010;R[27]=8'b0100_0110;
		R[28]=8'b0100_1010;R[29]=8'b0101_0010;R[30]=8'b0010_0010;
		R[31]=8'b0000_0000;R[32]=8'b0000_0000;//数字2
		
		R[33]=8'b0000_0000;R[34]=8'b0010_0010;R[35]=8'b0100_0001;
		R[36]=8'b0100_1001;R[37]=8'b0100_1001;R[38]=8'b0011_0110;
		R[39]=8'b0000_0000;R[40]=8'b0000_0000;//数字3
		
		R[41]=8'b0000_0100;R[42]=8'b0000_1100;R[43]=8'b0001_0100;
		R[44]=8'b0010_0100;R[45]=8'b0111_1111;R[46]=8'b0000_0100;
		R[47]=8'b0000_0000;R[48]=8'b0000_0000;//数字4

		R[49]=8'b0100_0010;R[50]=8'b0010_0100;R[51]=8'b0001_1000;
		R[52]=8'b0001_1000;R[53]=8'b0010_0100;R[54]=8'b0100_0010;
		R[55]=8'b1000_0001;R[56]=8'b0000_0000;//X
		
		r[97]=16'b1000_0000_0000_0001;//门开启
		r[98]=16'b1111_1111_1111_1111;//门关闭（全亮）
		r[99]=16'b0000_0000_0000_0000;R[99]=8'b0000_0000;//全灭
	end
	
always @(posedge clk2)//开关门动画和指示灯
begin
	r[15]={!Fin_4dn,!Fin_3up,!Fin_3dn,!Fin_2up,!Fin_2dn,!Fin_1up,4'b0000,!Fin_4,!Fin_3,!Fin_2,!Fin_1};//指示灯
	if (door==0)//如果需要开门，门逐渐打开
		case (cnt_d)
		2'b00:cnt_d<=2'b01;
		2'b01:cnt_d<=2'b10;
		2'b10:cnt_d<=2'b11;
		2'b11:cnt_d<=2'b11;
		default:cnt_d<=2'b11;
		endcase
	else 
		case (cnt_d)//如果需要开门，门逐渐关闭
		2'b00:cnt_d<=2'b00;
		2'b01:cnt_d<=2'b00;
		2'b10:cnt_d<=2'b01;
		2'b11:cnt_d<=2'b10;
		default:cnt_d<=2'b00;
		endcase
end

always @(posedge clk1)//根据状态对行寄存器进行赋值
begin
	begin
	if (err)//故障，显示X
	begin r[0][7:0]=R[49];r[1][7:0]=R[50];r[2][7:0]=R[51];r[3][7:0]=R[52];r[4][7:0]=R[53];r[5][7:0]=R[54];r[6][7:0]=R[55];end
	else
	case (drc)//运行方向，上行显示上箭头，下行显示下箭头，等待显示横杠
	2'b00:begin r[0][7:0]=R[16];r[1][7:0]=R[16];r[2][7:0]=R[16];r[3][7:0]=R[16];r[4][7:0]=R[16];r[5][7:0]=R[16];r[6][7:0]=R[99];end
	2'b01:begin r[0][7:0]=R[0];r[1][7:0]=R[1];r[2][7:0]=R[2];r[3][7:0]=R[3];r[4][7:0]=R[4];r[5][7:0]=R[5];r[6][7:0]=R[6];end
	2'b10:begin r[0][7:0]=R[8];r[1][7:0]=R[9];r[2][7:0]=R[10];r[3][7:0]=R[11];r[4][7:0]=R[12];r[5][7:0]=R[13];r[6][7:0]=R[14];end
	default:;
	endcase
	end
	case (c_floor)//当前楼层（1、2、3、4）
	2'b00:begin r[0][15:8]=R[17];r[1][15:8]=R[18];r[2][15:8]=R[19];r[3][15:8]=R[20];r[4][15:8]=R[21];r[5][15:8]=R[22];r[6][15:8]=R[23];end
	2'b01:begin r[0][15:8]=R[25];r[1][15:8]=R[26];r[2][15:8]=R[27];r[3][15:8]=R[28];r[4][15:8]=R[29];r[5][15:8]=R[30];r[6][15:8]=R[31];end
	2'b10:begin r[0][15:8]=R[33];r[1][15:8]=R[34];r[2][15:8]=R[35];r[3][15:8]=R[36];r[4][15:8]=R[37];r[5][15:8]=R[38];r[6][15:8]=R[39];end
	2'b11:begin r[0][15:8]=R[41];r[1][15:8]=R[42];r[2][15:8]=R[43];r[3][15:8]=R[44];r[4][15:8]=R[45];r[5][15:8]=R[46];r[6][15:8]=R[47];end
	default:;
	endcase
	case (cnt_d)//开关门的动画
	2'b00:begin r[7]=r[98]; r[8]=r[98]; r[9]=r[98]; r[10]=r[98]; r[11]=r[98]; r[12]=r[98]; r[13]=r[98]; r[14]=r[98];end
	2'b01:begin r[7]=r[98]; r[8]=r[98]; r[9]=r[98]; r[10]=r[97]; r[11]=r[97]; r[12]=r[98]; r[13]=r[98]; r[14]=r[98];end
	2'b10:begin r[7]=r[98]; r[8]=r[98]; r[9]=r[97]; r[10]=r[97]; r[11]=r[97]; r[12]=r[97]; r[13]=r[98]; r[14]=r[98];end
	2'b11:begin r[7]=r[98]; r[8]=r[97]; r[9]=r[97]; r[10]=r[97]; r[11]=r[97]; r[12]=r[97]; r[13]=r[97]; r[14]=r[98];end
	default:;
	endcase
end

always @(posedge clk1)//点阵扫描
	begin
	col<=col+1'b1;
	begin
	case(col)
	4'b0000:row=r[0];
	4'b0001:row=r[1];
	4'b0010:row=r[2];
	4'b0011:row=r[3];
	4'b0100:row=r[4];
	4'b0101:row=r[5];
	4'b0110:row=r[6];
	4'b0111:row=r[7];
	4'b1000:row=r[8];
	4'b1001:row=r[9];
	4'b1010:row=r[10];
	4'b1011:row=r[11];
	4'b1100:row=r[12];
	4'b1101:row=r[13];
	4'b1110:row=r[14];
	4'b1111:row=r[15];
	default:row=r[97];
	endcase
	end
	end


always @(posedge clk)//内部分频
begin
      if (i==10000/2-1)  
           begin
             i<=0; clk1<=~clk1;
           end
        else  i<=i+1;
end

always @(posedge clk)//内部分频
begin
        if (j==5000000/2-1)  
           begin
             j<=0; clk2<=~clk2;
           end
        else  j<=j+1;
end
endmodule
