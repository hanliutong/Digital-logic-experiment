library verilog;
use verilog.vl_types.all;
entity shifting_register_vlg_vec_tst is
end shifting_register_vlg_vec_tst;
