library verilog;
use verilog.vl_types.all;
entity keyboard_shake_vlg_vec_tst is
end keyboard_shake_vlg_vec_tst;
