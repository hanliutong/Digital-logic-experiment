library verilog;
use verilog.vl_types.all;
entity SEL6_vlg_vec_tst is
end SEL6_vlg_vec_tst;
