library verilog;
use verilog.vl_types.all;
entity project6_vlg_vec_tst is
end project6_vlg_vec_tst;
