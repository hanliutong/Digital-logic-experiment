library verilog;
use verilog.vl_types.all;
entity dynamic_scanning_vlg_vec_tst is
end dynamic_scanning_vlg_vec_tst;
