library verilog;
use verilog.vl_types.all;
entity decoder2_4_vlg_check_tst is
    port(
        out1            : in     vl_logic;
        out2            : in     vl_logic;
        out3            : in     vl_logic;
        out4            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder2_4_vlg_check_tst;
