library verilog;
use verilog.vl_types.all;
entity project7_vlg_vec_tst is
end project7_vlg_vec_tst;
